module comProc_tb();
	
endmodule